PACKAGE mydefinitions IS
    CONSTANT add : INTEGER := 0;
    CONSTANT subt : INTEGER := 1;
    CONSTANT neg : INTEGER := 2;
    CONSTANT mul : INTEGER := 3;
    CONSTANT div : INTEGER := 4;
    CONSTANT modu : INTEGER := 5;

    CONSTANT nicht : INTEGER := 6;
    CONSTANT und : INTEGER := 7;
    CONSTANT oder : INTEGER := 8;
    CONSTANT beq : INTEGER := 9;
    CONSTANT bneq : INTEGER := 10;
    CONSTANT blt : INTEGER := 11;
    CONSTANT jmp : INTEGER := 12;
    CONSTANT ldw : INTEGER := 13;
    CONSTANT stw : INTEGER := 14;

END PACKAGE mydefinitions;

