package mydefinitions is
    constant add : integer := 0;
    constant subt : integer := 1;
    constant neg : integer := 2;
    constant mul : integer := 3;
    constant div : integer := 4;
    constant modu : integer := 5;

    constant nicht : integer := 6;
    constant und : integer := 7;
    constant oder : integer := 8;
    constant beq : integer := 9;
    constant bneq : integer := 10;
    constant blt : integer := 11;
    constant jmp : integer := 12;
    constant ldw : integer := 13;
    constant stw : integer := 14;

end package mydefinitions;