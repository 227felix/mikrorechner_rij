package mydefinitions is
    constant add : integer := 0;
    constant subt : integer := 1;
    constant neg : integer := 2;

    constant nicht : integer := 3;
    constant und : integer := 4;
    constant oder : integer := 5;
    constant beq : integer := 6;
    constant bneq : integer := 7;
    constant blt : integer := 8;
    constant jmp : integer := 9;
    constant ldw : integer := 10;
    constant stw : integer := 11;
    constant mul : integer := 12;
    constant div : integer := 13;
    constant modu : integer := 14;

end package mydefinitions;